library verilog;
use verilog.vl_types.all;
entity Isaev11_vlg_vec_tst is
end Isaev11_vlg_vec_tst;
