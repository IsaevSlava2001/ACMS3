library verilog;
use verilog.vl_types.all;
entity Isaev12_vlg_vec_tst is
end Isaev12_vlg_vec_tst;
