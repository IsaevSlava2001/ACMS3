library verilog;
use verilog.vl_types.all;
entity Isaev21 is
    port(
        F               : out    vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        D0              : in     vl_logic;
        D2              : in     vl_logic;
        D1              : in     vl_logic;
        D3              : in     vl_logic;
        D5              : in     vl_logic;
        D4              : in     vl_logic;
        D6              : in     vl_logic;
        D7              : in     vl_logic
    );
end Isaev21;
