library verilog;
use verilog.vl_types.all;
entity Isaev23_vlg_vec_tst is
end Isaev23_vlg_vec_tst;
