library verilog;
use verilog.vl_types.all;
entity lab311_vlg_vec_tst is
end lab311_vlg_vec_tst;
