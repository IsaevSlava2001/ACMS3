library verilog;
use verilog.vl_types.all;
entity Isaev21_vlg_vec_tst is
end Isaev21_vlg_vec_tst;
