library verilog;
use verilog.vl_types.all;
entity Isaev22_vlg_vec_tst is
end Isaev22_vlg_vec_tst;
